module EXE_Stage(
    input clk, rst,
    input [31:0] pcIn,
    output [31:0] pc
);
endmodule