module IF_Stage(
    input clk, rst, freeze, branchTaken,
    input[31:0] branchAddress,
    output[31:0] pc, instruction);


endmodule