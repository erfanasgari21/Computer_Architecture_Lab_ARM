module EXE_Stage_Reg(
    input clk, rst,
    input [31:0] pcIn,
    output [31:0] pc
);

endmodule