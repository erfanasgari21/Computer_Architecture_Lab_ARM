module Val_Generator(
    input [31:0] valRm, shiftOperandImm
)